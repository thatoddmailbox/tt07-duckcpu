`default_nettype none

module spi(
	input wire clk,
	input wire rst
);

endmodule
